module test(a, b, output c);
input a;
input b;

wire w1;
wire w2;

and(c, a, b);

endmodule